`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Insituto Tecnol�gico de Costa Rica
// Students:
//  -Jose Antonio Espinoza Chaves 
//  -David Obando Pereira
//  -Rolando Vega Marino
//  -Naheem Johnson Sol�s
// Design Name: Sequential Multiplier
// Module Name: Shift register
//////////////////////////////////////////////////////////////////////////////////
module shiftRegister(clk, rst, Shift, load, Data_In, Data_Out);
    input clk, rst, Shift, load;
    input [3:0] Data_In;
    output reg [3:0] Data_Out;

always @(posedge clk or posedge rst)
    if (rst)
        Data_Out = 4'b0000;
    else if(Shift)
        Data_Out = {Data_Out[3], Data_Out[3:1]};
    else if(load)
        Data_Out = Data_In;
    else
        Data_Out = Data_Out;

endmodule